`timescale 1ns/1ps
`define DEF_LEAK 1
`define DEF_THRESHOLD 8

`define DEF_V_SIZE 3


/* 4-bit adder. 
 * valid input range: 0-15
 * If the result overflows, output will be 0b11111 meaning infinity
*/
module clipped_adder#(V_SIZE = `DEF_V_SIZE)(
    input unsigned [V_SIZE+1:0] a,
    input unsigned [V_SIZE+1:0] b,
    output unsigned [V_SIZE+1:0] out
);

wire unsigned [V_SIZE+1:0] sum;
assign sum = a + b;
assign out = a[V_SIZE+1] || b[V_SIZE+1] || sum[V_SIZE+1] ? {(V_SIZE+1){1'b1}} : sum;

endmodule

module lif_core#(V_SIZE = `DEF_V_SIZE)(
     input unsigned [V_SIZE:0] prev_v,
     input unsigned [V_SIZE+1:0] spike_in,
     input unsigned [V_SIZE:0] leak,
     output unsigned [V_SIZE+1:0] out
);

wire unsigned [V_SIZE+1:0] padded_v = {1'b0, prev_v};
wire unsigned [V_SIZE+1:0] padded_leak = {1'b0, leak};
wire unsigned [V_SIZE+1:0] sum;
wire unsigned [V_SIZE+1:0] ans;
assign sum = padded_v + spike_in;
assign ans = sum - padded_leak;

assign out = spike_in[V_SIZE+1] ? {(V_SIZE+1){1'b1}} : sum > padded_leak ?  ans[V_SIZE+1] ? {(V_SIZE+1){1'b1}} : ans : 0;

endmodule

module lif(V_SIZE = `DEF_V_SIZE, THRESHOLD = `DEF_THRESHOLD, LEAK = `DEF_LEAK)(
    input clk,
    input reset,
    input unsigned [V_SIZE+1:0] spike_in,
    output reg spike_out,
    output unsigned [V_SIZE:0] waveform
);

wire unsigned [V_SIZE+1:0] sum;
wire unsigned [V_SIZE:0] next_volt;
reg unsigned [V_SIZE:0] voltage;
wire has_spike;
wire unsigned [V_SIZE:0] leak = LEAK;
lif_core add(voltage, spike_in, leak, sum);
assign has_spike = sum >= THRESHOLD;
assign next_volt = has_spike ? 0 : sum;
assign waveform = voltage;

always @(posedge clk) begin
    if (reset) begin
        voltage <= 0;
        spike_out <= 0;
    end else begin
        voltage <= next_volt;
        spike_out <= has_spike;
    end
end

endmodule

module lif_sum3(V_SIZE = `DEF_V_SIZE, THRESHOLD = `DEF_THRESHOLD, LEAK = `DEF_LEAK)(
    input clk,
    input reset,
    input unsigned [V_SIZE+1:0] i1,
    input unsigned [V_SIZE+1:0] i2,
    input unsigned [V_SIZE+1:0] i3,
    output spike,
    output unsigned [V_SIZE+1:0] waveform
);

wire unsigned [V_SIZE+1:0] i12;
wire unsigned [V_SIZE+1:0] i123;
clipped_adder #(V_SIZE) a1(i1, i2, i12);
clipped_adder #(V_SIZE) a2(i12, i3, i123);
lif #(V_SIZE, THRESHOLD, LEAK) ni(clk, reset, i123, spike, waveform);

endmodule

module wrapper(
    input clk,
    input reset,
    input s1,
    input s2,
    input s3,
    output spike,
    output unsigned [`V_SIZE:0] waveform
);

wire unsigned [`I_SIZE:0] i1 = s1 ? `W1 : 0;
wire unsigned [`I_SIZE:0] i2 = s2 ? `W2 : 0;
wire unsigned [`I_SIZE:0] i3 = s3 ? `W3 : 0;
wire unsigned [`I_SIZE:0] i12;
wire unsigned [`I_SIZE:0] i123;

clipped_adder a1(i1, i2, i12);
clipped_adder a2(i12, i3, i123);

lif ni(clk, reset, i123, spike, waveform);

endmodule